logic [23:0] x_re [0:1023] = {    24'b111111111111011101110000,	//-0.000261
								   24'b111111111111101100010101,	//-0.000150 
								   24'b000000000000001000010101,	//0.000064 
								   24'b000000000000000110100101,	//0.000050 
								   24'b111111111111110101100110,	//-0.000079 
								   24'b111111111111111110100100,	//-0.000011 
								   24'b000000000000010011001101,	//0.000147 
								   24'b000000000000000001001111,	//0.000009 
								   24'b111111111111000101010001,	//-0.000448 
								   24'b111111111111111011000001,	//-0.000038 
								   24'b111111111110101010100010,	//-0.000652 
								   24'b111111111111000100001101,	//-0.000456 
								   24'b000000000000011110011001,	//0.000232 
								   24'b000000000000010000011100,	//0.000125 
								   24'b111111111110111100110101,	//-0.000512 
								   24'b111111111111100100000010,	//-0.000213 
								   24'b111111111111100010100100,	//-0.000225 
								   24'b000000000001001010011000,	//0.000567 
								   24'b111111111110100111011010,	//-0.000676 
								   24'b111111111101100100100101,	//-0.001186 
								   24'b000000000001000100011000,	//0.000522 
								   24'b111111111110010011110010,	//-0.000826 
								   24'b000000000000010111000111,	//0.000176 
								   24'b000000000000000010101110,	//0.000021 
								   24'b000000000000001100010001,	//0.000094 
								   24'b000000000000000011100000,	//0.000027 
								   24'b111111111111111110101000,	//-0.000010 
								   24'b000000000000010000011000,	//0.000125 
								   24'b111111111111111101111000,	//-0.000016 
								   24'b111111111111011111100110,	//-0.000247 
								   24'b000000000000100011100110,	//0.000272 
								   24'b000000000000000110101001,	//0.000051 
								   24'b111111111111111100100110,	//-0.000026 
								   24'b000000000000010001001001,	//0.000131 
								   24'b000000000000000010010000,	//0.000017 
								   24'b111111111111110100000011,	//-0.000091 
								   24'b000000000000000111101111,	//0.000059 
								   24'b000000000000000011011000,	//0.000026 
								   24'b000000000000011110001110,	//0.000231 
								   24'b111111111111110011100100,	//-0.000095 
								   24'b000000000000001010011001,	//0.000079 
								   24'b000000000000000010011001,	//0.000018 
								   24'b000000000000011001111001,	//0.000198 
								   24'b111111111111111110010011,	//-0.000013 
								   24'b111111111111111010111010,	//-0.000039 
								   24'b000000000000001001101101,	//0.000074 
								   24'b000000000000011001010011,	//0.000193 
								   24'b111111111111111110011001,	//-0.000012 
								   24'b111111111111110111110010,	//-0.000063 
								   24'b111111111111111110110100,	//-0.000009 
								   24'b000000000000000010110011,	//0.000021 
								   24'b111111111111111100110110,	//-0.000024 
								   24'b111111111111110111000101,	//-0.000068 
								   24'b000000000000001011011111,	//0.000088 
								   24'b000000000000011101001101,	//0.000223 
								   24'b111111111111110101101000,	//-0.000079 
								   24'b000000000000000011011101,	//0.000026 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111110000011010,	//-0.000119 
								   24'b000000000000010101000011,	//0.000161 
								   24'b000000000000011001101110,	//0.000196 
								   24'b000000000000000110000111,	//0.000047 
								   24'b111111111111101110011000,	//-0.000134 
								   24'b111111111111111100111000,	//-0.000024 
								   24'b111111111111111011101011,	//-0.000033 
								   24'b000000000000010101000111,	//0.000161 
								   24'b000000000000000000110101,	//0.000006 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b000000000000000011000010,	//0.000023 
								   24'b000000000000000011100101,	//0.000027 
								   24'b000000000000000000110111,	//0.000007 
								   24'b000000000000011110100001,	//0.000233 
								   24'b111111111111111001101011,	//-0.000048 
								   24'b000000000000000110110101,	//0.000052 
								   24'b000000000000000011100110,	//0.000027 
								   24'b111111111111100011100010,	//-0.000217 
								   24'b111111111111110111000011,	//-0.000068 
								   24'b111111111111110010110010,	//-0.000101 
								   24'b111111111111111100001011,	//-0.000029 
								   24'b111111111111110110010110,	//-0.000074 
								   24'b000000000000001000111111,	//0.000069 
								   24'b000000000000000100101101,	//0.000036 
								   24'b111111111111111100001011,	//-0.000029 
								   24'b111111111111111010111011,	//-0.000039 
								   24'b000000000000000110010100,	//0.000048 
								   24'b000000000000000000010011,	//0.000002 
								   24'b000000000000000001000101,	//0.000008 
								   24'b000000000000000001110011,	//0.000014 
								   24'b000000000000010110001001,	//0.000169 
								   24'b000000000000010001101010,	//0.000135 
								   24'b000000000000001010010100,	//0.000079 
								   24'b111111111111011111101100,	//-0.000247 
								   24'b111111111111110111101111,	//-0.000063 
								   24'b000000000000001011101000,	//0.000089 
								   24'b111111111111101100111100,	//-0.000145 
								   24'b000000000000001010100111,	//0.000081 
								   24'b000000000000000010011001,	//0.000018 
								   24'b111111111111111001000010,	//-0.000053 
								   24'b000000000000001110001111,	//0.000109 
								   24'b000000000000001000101110,	//0.000067 
								   24'b111111111111110110011010,	//-0.000073 
								   24'b000000000000000110001000,	//0.000047 
								   24'b111111111111110111000001,	//-0.000069 
								   24'b000000000000000001100001,	//0.000012 
								   24'b111111111111111110100101,	//-0.000011 
								   24'b111111111111111101011111,	//-0.000019 
								   24'b111111111111111110001110,	//-0.000014 
								   24'b111111111111111110001000,	//-0.000014 
								   24'b111111111111111101111010,	//-0.000016 
								   24'b111111111111111101111111,	//-0.000015 
								   24'b111111111111111110000000,	//-0.000015 
								   24'b000000000000000000010110,	//0.000003 
								   24'b000000000000000000101011,	//0.000005 
								   24'b111111111111111111000011,	//-0.000007 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b000000000000000010110111,	//0.000022 
								   24'b000000000000000000110110,	//0.000006 
								   24'b111111111111111101001001,	//-0.000022 
								   24'b111111111111111110101001,	//-0.000010 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000010010000,	//0.000017 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b111111111111111101000000,	//-0.000023 
								   24'b000000000000000001100101,	//0.000012 
								   24'b000000000000000001111010,	//0.000015 
								   24'b000000000000000000001011,	//0.000001 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111101001110,	//-0.000021 
								   24'b000000000000000000110010,	//0.000006 
								   24'b000000000000000001000011,	//0.000008 
								   24'b000000000000000000001101,	//0.000002 
								   24'b000000000000000000111101,	//0.000007 
								   24'b000000000000000000000001,	//0.000000 
								   24'b000000000000000000000110,	//0.000001 
								   24'b000000000000000001110111,	//0.000014 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111110000011,	//-0.000015 
								   24'b000000000000000010011011,	//0.000018 
								   24'b000000000000000000110011,	//0.000006 
								   24'b000000000000000010000111,	//0.000016 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b000000000000000000000010,	//0.000000 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b000000000000000000011111,	//0.000004 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b000000000000000000010011,	//0.000002 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b000000000000000000000000,	//-0.000000 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000100111,	//0.000005 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111110101010,	//-0.000010 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b000000000000000000110101,	//0.000006 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b000000000000000000001101,	//0.000001 
								   24'b000000000000000000010001,	//0.000002 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111011010,	//-0.000005 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b000000000000000000011011,	//0.000003 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000101011,	//0.000005 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b000000000000000000010000,	//0.000002 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000000011,	//0.000000 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000011100,	//0.000003 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b000000000000000000001100,	//0.000001 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b000000000000000000001110,	//0.000002 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111100011,	//-0.000004 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111011010,	//-0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b000000000000000000000100,	//0.000000 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111110111101,	//-0.000008 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b000000000000000000010110,	//0.000003 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000000111,	//0.000001 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111000011,	//-0.000007 
								   24'b000000000000000000000010,	//0.000000 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b000000000000000000010001,	//0.000002 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b000000000000000000010111,	//0.000003 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b000000000000000000000001,	//0.000000 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b000000000000000000000001,	//0.000000 
								   24'b000000000000000000001000,	//0.000001 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111110111001,	//-0.000008 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111110101011,	//-0.000010 
								   24'b000000000000000000111111,	//0.000008 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b000000000000000000011011,	//0.000003 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b000000000000000000101001,	//0.000005 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b000000000000000000001000,	//0.000001 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b000000000000000001001011,	//0.000009 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b000000000000000000100100,	//0.000004 
								   24'b111111111111111110111011,	//-0.000008 
								   24'b111111111111111110011101,	//-0.000012 
								   24'b000000000000000000110011,	//0.000006 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b111111111111111110110000,	//-0.000010 
								   24'b000000000000000000101000,	//0.000005 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000000001010,	//0.000001 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b000000000000000001100011,	//0.000012 
								   24'b000000000000000000011011,	//0.000003 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b000000000000000000010010,	//0.000002 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b000000000000000000111111,	//0.000008 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000000010,	//0.000000 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b000000000000000000100010,	//0.000004 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b000000000000000001001100,	//0.000009 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111110111010,	//-0.000008 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111110110010,	//-0.000009 
								   24'b000000000000000000111110,	//0.000007 
								   24'b111111111111111110110010,	//-0.000009 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111110111010,	//-0.000008 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b000000000000000001001100,	//0.000009 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b000000000000000000100010,	//0.000004 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b000000000000000000000010,	//0.000000 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000101000,	//0.000005 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b000000000000000000111111,	//0.000008 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b000000000000000000010010,	//0.000002 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000010100,	//0.000002 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000001100011,	//0.000012 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b000000000000000000001010,	//0.000001 
								   24'b000000000000000000010000,	//0.000002 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b000000000000000000101000,	//0.000005 
								   24'b111111111111111110110000,	//-0.000010 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b000000000000000000110011,	//0.000006 
								   24'b111111111111111110011101,	//-0.000012 
								   24'b111111111111111110111011,	//-0.000008 
								   24'b000000000000000000100100,	//0.000004 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b000000000000000001001011,	//0.000009 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b000000000000000000001000,	//0.000001 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b000000000000000000101001,	//0.000005 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b000000000000000000011011,	//0.000003 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b000000000000000000111111,	//0.000008 
								   24'b111111111111111110101011,	//-0.000010 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111110111001,	//-0.000008 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b000000000000000000001000,	//0.000001 
								   24'b000000000000000000000001,	//0.000000 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b000000000000000000000000,	//0.000000 
								   24'b000000000000000000000001,	//0.000000 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b000000000000000000010111,	//0.000003 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b000000000000000000010001,	//0.000002 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b000000000000000000000010,	//0.000000 
								   24'b111111111111111111000011,	//-0.000007 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b000000000000000000000111,	//0.000001 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b000000000000000000010110,	//0.000003 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111110111101,	//-0.000008 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b000000000000000000000100,	//0.000000 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111011010,	//-0.000004 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111100011,	//-0.000004 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b000000000000000000001110,	//0.000002 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b000000000000000000001100,	//0.000001 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b000000000000000000011100,	//0.000003 
								   24'b000000000000000000010100,	//0.000002 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b000000000000000000000011,	//0.000000 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b000000000000000000010000,	//0.000002 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b000000000000000000101011,	//0.000005 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b000000000000000000011011,	//0.000003 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111011010,	//-0.000005 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000001101,	//0.000001 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000110101,	//0.000006 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111110101010,	//-0.000010 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b000000000000000000100111,	//0.000005 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b000000000000000000000000,	//-0.000000 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b000000000000000000010011,	//0.000002 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b000000000000000000011111,	//0.000004 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b000000000000000000000010,	//0.000000 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b000000000000000010000111,	//0.000016 
								   24'b000000000000000000110011,	//0.000006 
								   24'b000000000000000010011011,	//0.000018 
								   24'b111111111111111110000011,	//-0.000015 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b000000000000000001110111,	//0.000014 
								   24'b000000000000000000000110,	//0.000001 
								   24'b000000000000000000000001,	//0.000000 
								   24'b000000000000000000111101,	//0.000007 
								   24'b000000000000000000001101,	//0.000002 
								   24'b000000000000000001000011,	//0.000008 
								   24'b000000000000000000110010,	//0.000006 
								   24'b111111111111111101001110,	//-0.000021 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b000000000000000000001011,	//0.000001 
								   24'b000000000000000001111010,	//0.000015 
								   24'b000000000000000001100101,	//0.000012 
								   24'b111111111111111101000000,	//-0.000023 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b000000000000000010010000,	//0.000017 
								   24'b000000000000000000011011,	//0.000003 
								   24'b111111111111111110101001,	//-0.000010 
								   24'b111111111111111101001001,	//-0.000022 
								   24'b000000000000000000110110,	//0.000006 
								   24'b000000000000000010110111,	//0.000022 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111000011,	//-0.000007 
								   24'b000000000000000000101011,	//0.000005 
								   24'b000000000000000000010110,	//0.000003 
								   24'b111111111111111110000000,	//-0.000015 
								   24'b111111111111111101111111,	//-0.000015 
								   24'b111111111111111101111010,	//-0.000016 
								   24'b111111111111111110001000,	//-0.000014 
								   24'b111111111111111110001110,	//-0.000014 
								   24'b111111111111111101011111,	//-0.000019 
								   24'b111111111111111110100101,	//-0.000011 
								   24'b000000000000000001100001,	//0.000012 
								   24'b111111111111110111000001,	//-0.000069 
								   24'b000000000000000110001000,	//0.000047 
								   24'b111111111111110110011010,	//-0.000073 
								   24'b000000000000001000101110,	//0.000067 
								   24'b000000000000001110001111,	//0.000109 
								   24'b111111111111111001000010,	//-0.000053 
								   24'b000000000000000010011001,	//0.000018 
								   24'b000000000000001010100111,	//0.000081 
								   24'b111111111111101100111100,	//-0.000145 
								   24'b000000000000001011101000,	//0.000089 
								   24'b111111111111110111101111,	//-0.000063 
								   24'b111111111111011111101100,	//-0.000247 
								   24'b000000000000001010010100,	//0.000079 
								   24'b000000000000010001101010,	//0.000135 
								   24'b000000000000010110001001,	//0.000169 
								   24'b000000000000000001110011,	//0.000014 
								   24'b000000000000000001000101,	//0.000008 
								   24'b000000000000000000010011,	//0.000002 
								   24'b000000000000000110010100,	//0.000048 
								   24'b111111111111111010111011,	//-0.000039 
								   24'b111111111111111100001011,	//-0.000029 
								   24'b000000000000000100101101,	//0.000036 
								   24'b000000000000001000111111,	//0.000069 
								   24'b111111111111110110010110,	//-0.000074 
								   24'b111111111111111100001011,	//-0.000029 
								   24'b111111111111110010110010,	//-0.000101 
								   24'b111111111111110111000011,	//-0.000068 
								   24'b111111111111100011100010,	//-0.000217 
								   24'b000000000000000011100110,	//0.000027 
								   24'b000000000000000110110101,	//0.000052 
								   24'b111111111111111001101011,	//-0.000048 
								   24'b000000000000011110100001,	//0.000233 
								   24'b000000000000000000110111,	//0.000007 
								   24'b000000000000000011100101,	//0.000027 
								   24'b000000000000000011000010,	//0.000023 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b000000000000000000110101,	//0.000006 
								   24'b000000000000010101000111,	//0.000161 
								   24'b111111111111111011101011,	//-0.000033 
								   24'b111111111111111100111000,	//-0.000024 
								   24'b111111111111101110011000,	//-0.000134 
								   24'b000000000000000110000111,	//0.000047 
								   24'b000000000000011001101110,	//0.000196 
								   24'b000000000000010101000011,	//0.000161 
								   24'b111111111111110000011010,	//-0.000119 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b000000000000000011011101,	//0.000026 
								   24'b111111111111110101101000,	//-0.000079 
								   24'b000000000000011101001101,	//0.000223 
								   24'b000000000000001011011111,	//0.000088 
								   24'b111111111111110111000101,	//-0.000068 
								   24'b111111111111111100110110,	//-0.000024 
								   24'b000000000000000010110011,	//0.000021 
								   24'b111111111111111110110100,	//-0.000009 
								   24'b111111111111110111110010,	//-0.000063 
								   24'b111111111111111110011001,	//-0.000012 
								   24'b000000000000011001010011,	//0.000193 
								   24'b000000000000001001101101,	//0.000074 
								   24'b111111111111111010111010,	//-0.000039 
								   24'b111111111111111110010011,	//-0.000013 
								   24'b000000000000011001111001,	//0.000198 
								   24'b000000000000000010011001,	//0.000018 
								   24'b000000000000001010011001,	//0.000079 
								   24'b111111111111110011100100,	//-0.000095 
								   24'b000000000000011110001110,	//0.000231 
								   24'b000000000000000011011000,	//0.000026 
								   24'b000000000000000111101111,	//0.000059 
								   24'b111111111111110100000011,	//-0.000091 
								   24'b000000000000000010010000,	//0.000017 
								   24'b000000000000010001001001,	//0.000131 
								   24'b111111111111111100100110,	//-0.000026 
								   24'b000000000000000110101001,	//0.000051 
								   24'b000000000000100011100110,	//0.000272 
								   24'b111111111111011111100110,	//-0.000247 
								   24'b111111111111111101111000,	//-0.000016 
								   24'b000000000000010000011000,	//0.000125 
								   24'b111111111111111110101000,	//-0.000010 
								   24'b000000000000000011100000,	//0.000027 
								   24'b000000000000001100010001,	//0.000094 
								   24'b000000000000000010101110,	//0.000021 
								   24'b000000000000010111000111,	//0.000176 
								   24'b111111111110010011110010,	//-0.000826 
								   24'b000000000001000100011000,	//0.000522 
								   24'b111111111101100100100101,	//-0.001186 
								   24'b111111111110100111011010,	//-0.000676 
								   24'b000000000001001010011000,	//0.000567 
								   24'b111111111111100010100100,	//-0.000225 
								   24'b111111111111100100000010,	//-0.000213 
								   24'b111111111110111100110101,	//-0.000512 
								   24'b000000000000010000011100,	//0.000125 
								   24'b000000000000011110011001,	//0.000232 
								   24'b111111111111000100001101,	//-0.000456 
								   24'b111111111110101010100010,	//-0.000652 
								   24'b111111111111111011000001,	//-0.000038 
								   24'b111111111111000101010001,	//-0.000448 
								   24'b000000000000000001001111,	//0.000009 
								   24'b000000000000010011001101,	//0.000147 
								   24'b111111111111111110100100,	//-0.000011 
								   24'b111111111111110101100110,	//-0.000079 
								   24'b000000000000000110100101,	//0.000050 
								   24'b000000000000001000010101,	//0.000064 
								   24'b111111111111101100010101};	//-0.000150 


logic [23:0] x_im [0:1023] = {     24'b000000000000000000000000,	//0.000000
								   24'b000000000000000001101100,	//0.000013 
								   24'b000000000000000010011011,	//0.000019 
								   24'b000000000000000010000010,	//0.000015 
								   24'b111111111111110101001001,	//-0.000083 
								   24'b000000000000000011100001,	//0.000027 
								   24'b111111111111110011011111,	//-0.000096 
								   24'b111111111111110110011100,	//-0.000073 
								   24'b111111111111011001101101,	//-0.000292 
								   24'b000000000000000001111111,	//0.000015 
								   24'b000000000001000101111111,	//0.000534 
								   24'b000000000000000010011111,	//0.000019 
								   24'b000000000000001000001001,	//0.000062 
								   24'b111111111110111100000011,	//-0.000518 
								   24'b000000000011000011010000,	//0.001490 
								   24'b111111111100100111100111,	//-0.001651 
								   24'b000000000011010111001100,	//0.001642 
								   24'b000000000000110111001101,	//0.000421 
								   24'b000000000000100100100001,	//0.000279 
								   24'b000000000000001010110110,	//0.000083 
								   24'b000000000000001111100110,	//0.000119 
								   24'b111111111110110011110000,	//-0.000582 
								   24'b111111111111100011111000,	//-0.000215 
								   24'b111111111111111011010101,	//-0.000036 
								   24'b000000000000000100000011,	//0.000031 
								   24'b000000000000001011110010,	//0.000090 
								   24'b111111111111111011101111,	//-0.000033 
								   24'b111111111111111110011001,	//-0.000012 
								   24'b111111111111110100111001,	//-0.000085 
								   24'b000000000000000100011111,	//0.000034 
								   24'b000000000001000110111000,	//0.000541 
								   24'b111111111111100101111010,	//-0.000199 
								   24'b111111111111100110001110,	//-0.000197 
								   24'b000000000000000110011010,	//0.000049 
								   24'b000000000000000110111110,	//0.000053 
								   24'b111111111111110110001110,	//-0.000075 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000001010010,	//0.000010 
								   24'b111111111111101110100011,	//-0.000133 
								   24'b000000000000001001000010,	//0.000069 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111101010101100,	//-0.000163 
								   24'b000000000000000010100110,	//0.000020 
								   24'b111111111111110111000110,	//-0.000068 
								   24'b111111111111111000100010,	//-0.000057 
								   24'b111111111111110011011011,	//-0.000096 
								   24'b111111111111010111101000,	//-0.000308 
								   24'b000000000000110011111100,	//0.000396 
								   24'b000000000000000111011110,	//0.000057 
								   24'b000000000000000111111111,	//0.000061 
								   24'b000000000000001110101001,	//0.000112 
								   24'b111111111111111101010101,	//-0.000020 
								   24'b000000000000001110111000,	//0.000113 
								   24'b000000000000000111110110,	//0.000060 
								   24'b000000000000001100111010,	//0.000098 
								   24'b111111111111111110101110,	//-0.000010 
								   24'b111111111111111110111000,	//-0.000009 
								   24'b111111111111110011101011,	//-0.000094 
								   24'b000000000000010010110100,	//0.000144 
								   24'b111111111111101011001011,	//-0.000159 
								   24'b111111111111101110110110,	//-0.000131 
								   24'b111111111111110100110010,	//-0.000086 
								   24'b111111111111111110001100,	//-0.000014 
								   24'b000000000000000111110110,	//0.000060 
								   24'b000000000000000000001110,	//0.000002 
								   24'b000000000000001000010110,	//0.000064 
								   24'b000000000000001010101111,	//0.000082 
								   24'b000000000000000101000000,	//0.000038 
								   24'b000000000000000000001011,	//0.000001 
								   24'b000000000000001010111001,	//0.000083 
								   24'b111111111111111010010000,	//-0.000044 
								   24'b111111111111110001010010,	//-0.000112 
								   24'b111111111111101110101000,	//-0.000133 
								   24'b000000000000001101010000,	//0.000101 
								   24'b000000000000011000111000,	//0.000190 
								   24'b111111111111110000010010,	//-0.000120 
								   24'b111111111111110010101100,	//-0.000102 
								   24'b111111111111111000000011,	//-0.000061 
								   24'b000000000000000010110101,	//0.000022 
								   24'b111111111111001110100111,	//-0.000377 
								   24'b111111111111111010001001,	//-0.000045 
								   24'b000000000000000010000101,	//0.000016 
								   24'b000000000000000100101110,	//0.000036 
								   24'b000000000000000100101111,	//0.000036 
								   24'b000000000000000010001000,	//0.000016 
								   24'b111111111111110001010110,	//-0.000112 
								   24'b111111111111111100100011,	//-0.000026 
								   24'b111111111111111010011110,	//-0.000042 
								   24'b000000000000001011111010,	//0.000091 
								   24'b000000000000010001011110,	//0.000133 
								   24'b000000000000001001001111,	//0.000070 
								   24'b000000000000000110011011,	//0.000049 
								   24'b000000000000000000000010,	//0.000000 
								   24'b000000000000000010100010,	//0.000019 
								   24'b111111111111110110101000,	//-0.000072 
								   24'b000000000000000001010101,	//0.000010 
								   24'b000000000000000101001111,	//0.000040 
								   24'b000000000000000000010000,	//0.000002 
								   24'b111111111111111001000000,	//-0.000053 
								   24'b000000000000001000110110,	//0.000067 
								   24'b000000000000000100111110,	//0.000038 
								   24'b000000000000001010111010,	//0.000083 
								   24'b000000000000000000110111,	//0.000007 
								   24'b111111111111111011001011,	//-0.000037 
								   24'b000000000000000101000011,	//0.000038 
								   24'b000000000000000011101111,	//0.000029 
								   24'b000000000000000100010110,	//0.000033 
								   24'b000000000000000010001111,	//0.000017 
								   24'b000000000000000010100000,	//0.000019 
								   24'b000000000000000100101100,	//0.000036 
								   24'b000000000000000110000110,	//0.000046 
								   24'b000000000000000110000000,	//0.000046 
								   24'b111111111111110111001100,	//-0.000067 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000001011,	//0.000001 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b000000000000001000010100,	//0.000063 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b000000000000000001011100,	//0.000011 
								   24'b000000000000000011001001,	//0.000024 
								   24'b111111111111111110101101,	//-0.000010 
								   24'b111111111111111101111111,	//-0.000015 
								   24'b000000000000000001001111,	//0.000009 
								   24'b000000000000000011000001,	//0.000023 
								   24'b000000000000000001010111,	//0.000010 
								   24'b000000000000000001101111,	//0.000013 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b000000000000000010100111,	//0.000020 
								   24'b111111111111111100110010,	//-0.000025 
								   24'b000000000000000010000001,	//0.000015 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b000000000000000010000100,	//0.000016 
								   24'b000000000000000010101001,	//0.000020 
								   24'b000000000000000010011101,	//0.000019 
								   24'b000000000000000001100000,	//0.000011 
								   24'b000000000000000000110001,	//0.000006 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b000000000000000010101011,	//0.000020 
								   24'b000000000000000010000010,	//0.000016 
								   24'b000000000000000001101110,	//0.000013 
								   24'b000000000000000001010000,	//0.000010 
								   24'b000000000000000001100001,	//0.000012 
								   24'b000000000000000001011000,	//0.000011 
								   24'b000000000000000010001000,	//0.000016 
								   24'b000000000000000001111000,	//0.000014 
								   24'b000000000000000001000001,	//0.000008 
								   24'b000000000000000001111100,	//0.000015 
								   24'b000000000000000001101001,	//0.000012 
								   24'b000000000000000001110001,	//0.000013 
								   24'b000000000000000001110010,	//0.000014 
								   24'b000000000000000001111011,	//0.000015 
								   24'b000000000000000000000111,	//0.000001 
								   24'b000000000000000000100100,	//0.000004 
								   24'b000000000000000001000011,	//0.000008 
								   24'b000000000000000000100111,	//0.000005 
								   24'b000000000000000001101010,	//0.000013 
								   24'b000000000000000000111001,	//0.000007 
								   24'b000000000000000000011101,	//0.000003 
								   24'b000000000000000001100000,	//0.000011 
								   24'b000000000000000001001011,	//0.000009 
								   24'b000000000000000001011110,	//0.000011 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000001011011,	//0.000011 
								   24'b000000000000000010000000,	//0.000015 
								   24'b000000000000000001101111,	//0.000013 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000111111,	//0.000008 
								   24'b000000000000000001000010,	//0.000008 
								   24'b000000000000000001001100,	//0.000009 
								   24'b000000000000000001000111,	//0.000008 
								   24'b000000000000000000111101,	//0.000007 
								   24'b000000000000000001010001,	//0.000010 
								   24'b000000000000000001001001,	//0.000009 
								   24'b000000000000000000111001,	//0.000007 
								   24'b000000000000000000111110,	//0.000007 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000001001010,	//0.000009 
								   24'b000000000000000000110110,	//0.000006 
								   24'b000000000000000001001001,	//0.000009 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000001000101,	//0.000008 
								   24'b000000000000000000001101,	//0.000001 
								   24'b000000000000000000100010,	//0.000004 
								   24'b000000000000000000110001,	//0.000006 
								   24'b000000000000000000110011,	//0.000006 
								   24'b000000000000000001001100,	//0.000009 
								   24'b000000000000000001100011,	//0.000012 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b000000000000000001001010,	//0.000009 
								   24'b000000000000000001001111,	//0.000009 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000110101,	//0.000006 
								   24'b000000000000000000110010,	//0.000006 
								   24'b000000000000000000111110,	//0.000007 
								   24'b000000000000000001001011,	//0.000009 
								   24'b000000000000000000100011,	//0.000004 
								   24'b000000000000000000110110,	//0.000006 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000001001111,	//0.000009 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000111100,	//0.000007 
								   24'b000000000000000000011100,	//0.000003 
								   24'b000000000000000000101111,	//0.000006 
								   24'b000000000000000001000000,	//0.000008 
								   24'b000000000000000000110100,	//0.000006 
								   24'b000000000000000001000001,	//0.000008 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000110110,	//0.000006 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000001001001,	//0.000009 
								   24'b000000000000000000010011,	//0.000002 
								   24'b000000000000000000101100,	//0.000005 
								   24'b000000000000000000110010,	//0.000006 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000111110,	//0.000007 
								   24'b000000000000000000100011,	//0.000004 
								   24'b000000000000000000110111,	//0.000007 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000111011,	//0.000007 
								   24'b000000000000000000100010,	//0.000004 
								   24'b000000000000000001001011,	//0.000009 
								   24'b000000000000000000010111,	//0.000003 
								   24'b000000000000000001000101,	//0.000008 
								   24'b000000000000000000110000,	//0.000006 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000000111110,	//0.000007 
								   24'b000000000000000000110011,	//0.000006 
								   24'b000000000000000000101100,	//0.000005 
								   24'b000000000000000000101100,	//0.000005 
								   24'b000000000000000000110010,	//0.000006 
								   24'b000000000000000000010110,	//0.000003 
								   24'b000000000000000000100111,	//0.000005 
								   24'b000000000000000000011101,	//0.000003 
								   24'b000000000000000000110111,	//0.000007 
								   24'b000000000000000000111011,	//0.000007 
								   24'b000000000000000000001111,	//0.000002 
								   24'b000000000000000000110110,	//0.000006 
								   24'b000000000000000000011000,	//0.000003 
								   24'b000000000000000000111010,	//0.000007 
								   24'b000000000000000000101110,	//0.000005 
								   24'b000000000000000000110000,	//0.000006 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000000101011,	//0.000005 
								   24'b000000000000000000110011,	//0.000006 
								   24'b000000000000000000101100,	//0.000005 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000001111,	//0.000002 
								   24'b000000000000000001000010,	//0.000008 
								   24'b000000000000000000001100,	//0.000001 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000100010,	//0.000004 
								   24'b000000000000000000110010,	//0.000006 
								   24'b000000000000000000111100,	//0.000007 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000100110,	//0.000005 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000000110100,	//0.000006 
								   24'b000000000000000000011100,	//0.000003 
								   24'b000000000000000000101111,	//0.000006 
								   24'b000000000000000000010011,	//0.000002 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000010110,	//0.000003 
								   24'b000000000000000000100100,	//0.000004 
								   24'b000000000000000000111101,	//0.000007 
								   24'b000000000000000000001101,	//0.000002 
								   24'b000000000000000000110110,	//0.000006 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000101111,	//0.000006 
								   24'b000000000000000000010111,	//0.000003 
								   24'b000000000000000000111010,	//0.000007 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000101111,	//0.000006 
								   24'b000000000000000000111100,	//0.000007 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000010101,	//0.000003 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000110111,	//0.000007 
								   24'b000000000000000000110100,	//0.000006 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000111000,	//0.000007 
								   24'b000000000000000000100101,	//0.000004 
								   24'b000000000000000000101101,	//0.000005 
								   24'b000000000000000000010111,	//0.000003 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000100101,	//0.000004 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000101011,	//0.000005 
								   24'b000000000000000000100100,	//0.000004 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000010101,	//0.000003 
								   24'b000000000000000000010101,	//0.000003 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000000010111,	//0.000003 
								   24'b000000000000000000110101,	//0.000006 
								   24'b000000000000000000001100,	//0.000001 
								   24'b000000000000000000111010,	//0.000007 
								   24'b000000000000000000011100,	//0.000003 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000000010101,	//0.000002 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000000100000,	//0.000004 
								   24'b000000000000000000001111,	//0.000002 
								   24'b000000000000000000101000,	//0.000005 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000000010110,	//0.000003 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000110000,	//0.000006 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000011010,	//0.000003 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000100011,	//0.000004 
								   24'b000000000000000000110000,	//0.000006 
								   24'b000000000000000000010011,	//0.000002 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000011000,	//0.000003 
								   24'b000000000000000000100000,	//0.000004 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000100111,	//0.000005 
								   24'b000000000000000000100100,	//0.000004 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000010101,	//0.000002 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000010010,	//0.000002 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000100101,	//0.000004 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000110001,	//0.000006 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000001011,	//0.000001 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b000000000000000000011000,	//0.000003 
								   24'b000000000000000000100011,	//0.000004 
								   24'b000000000000000000010111,	//0.000003 
								   24'b000000000000000000101010,	//0.000005 
								   24'b000000000000000000010110,	//0.000003 
								   24'b000000000000000000011100,	//0.000003 
								   24'b000000000000000000000111,	//0.000001 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000010101,	//0.000003 
								   24'b000000000000000000010010,	//0.000002 
								   24'b000000000000000000100000,	//0.000004 
								   24'b000000000000000000001011,	//0.000001 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000001110,	//0.000002 
								   24'b000000000000000000001000,	//0.000001 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000010101,	//0.000002 
								   24'b000000000000000000100011,	//0.000004 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000001010,	//0.000001 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000000010,	//0.000000 
								   24'b000000000000000000011010,	//0.000003 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000100100,	//0.000004 
								   24'b000000000000000000011000,	//0.000003 
								   24'b000000000000000000011110,	//0.000004 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b000000000000000000010010,	//0.000002 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000001110,	//0.000002 
								   24'b000000000000000000001111,	//0.000002 
								   24'b000000000000000000101111,	//0.000006 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000010101,	//0.000002 
								   24'b000000000000000000100010,	//0.000004 
								   24'b000000000000000000100010,	//0.000004 
								   24'b000000000000000000011111,	//0.000004 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000110011,	//0.000006 
								   24'b000000000000000000000100,	//0.000000 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b000000000000000000001010,	//0.000001 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000100101,	//0.000004 
								   24'b000000000000000000000100,	//0.000000 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b000000000000000000001010,	//0.000001 
								   24'b000000000000000000000110,	//0.000001 
								   24'b000000000000000000111011,	//0.000007 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000011001,	//0.000003 
								   24'b000000000000000000100110,	//0.000004 
								   24'b000000000000000000100101,	//0.000004 
								   24'b000000000000000000111010,	//0.000007 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000001011,	//0.000001 
								   24'b000000000000000000001000,	//0.000001 
								   24'b000000000000000000010101,	//0.000003 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b000000000000000000000111,	//0.000001 
								   24'b000000000000000000000000,	//-0.000000 
								   24'b000000000000000000111110,	//0.000007 
								   24'b000000000000000000011011,	//0.000003 
								   24'b000000000000000000010110,	//0.000003 
								   24'b000000000000000001001010,	//0.000009 
								   24'b000000000000000000010010,	//0.000002 
								   24'b000000000000000000100100,	//0.000004 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000000011,	//0.000000 
								   24'b000000000000000000101101,	//0.000005 
								   24'b111111111111111111011010,	//-0.000005 
								   24'b000000000000000000000100,	//0.000000 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111011010,	//-0.000005 
								   24'b000000000000000000011101,	//0.000003 
								   24'b000000000000000000110000,	//0.000006 
								   24'b000000000000000000010011,	//0.000002 
								   24'b000000000000000000001011,	//0.000001 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000110100,	//0.000006 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000111001,	//0.000007 
								   24'b000000000000000000000010,	//0.000000 
								   24'b000000000000000000101101,	//0.000005 
								   24'b000000000000000000100111,	//0.000005 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b000000000000000000101111,	//0.000006 
								   24'b000000000000000000011111,	//0.000004 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b000000000000000000101001,	//0.000005 
								   24'b000000000000000000001010,	//0.000001 
								   24'b000000000000000000001010,	//0.000001 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111011101,	//-0.000004 
								   24'b000000000000000000011010,	//0.000003 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b000000000000000000001101,	//0.000002 
								   24'b000000000000000000110100,	//0.000006 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b000000000000000000011000,	//0.000003 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b000000000000000000110010,	//0.000006 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b000000000000000000010011,	//0.000002 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b000000000000000000001001,	//0.000001 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b000000000000000000101110,	//0.000005 
								   24'b000000000000000000010100,	//0.000002 
								   24'b111111111111111111111111,	//-0.000000 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b000000000000000000100101,	//0.000004 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b000000000000000000010001,	//0.000002 
								   24'b000000000000000000011010,	//0.000003 
								   24'b000000000000000000101110,	//0.000005 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000001100,	//0.000001 
								   24'b000000000000000000110000,	//0.000006 
								   24'b000000000000000000101101,	//0.000005 
								   24'b000000000000000001001101,	//0.000009 
								   24'b000000000000000000100001,	//0.000004 
								   24'b000000000000000000000000,	//-0.000000 
								   24'b000000000000000000010101,	//0.000003 
								   24'b000000000000000000000111,	//0.000001 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b000000000000000000111000,	//0.000007 
								   24'b000000000000000000111010,	//0.000007 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b000000000000000000000010,	//0.000000 
								   24'b000000000000000000000110,	//0.000001 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b000000000000000000101011,	//0.000005 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b000000000000000000001101,	//0.000002 
								   24'b000000000000000000011000,	//0.000003 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111100011,	//-0.000004 
								   24'b000000000000000001000000,	//0.000008 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000001001,	//0.000001 
								   24'b000000000000000000001101,	//0.000002 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b000000000000000000001111,	//0.000002 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b000000000000000000101110,	//0.000005 
								   24'b000000000000000000010000,	//0.000002 
								   24'b000000000000000000010010,	//0.000002 
								   24'b000000000000000000110010,	//0.000006 
								   24'b000000000000000000100000,	//0.000004 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b000000000000000000011110,	//0.000004 
								   24'b000000000000000000100000,	//0.000004 
								   24'b000000000000000000111001,	//0.000007 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b000000000000000000010101,	//0.000003 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b000000000000000001000000,	//0.000008 
								   24'b000000000000000000101000,	//0.000005 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b000000000000000000001100,	//0.000001 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000001001,	//0.000001 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b000000000000000000011101,	//0.000004 
								   24'b000000000000000000001100,	//0.000001 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b000000000000000000110000,	//0.000006 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b000000000000000000100001,	//0.000004 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b000000000000000000010000,	//0.000002 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b000000000000000000000101,	//0.000001 
								   24'b000000000000000000011110,	//0.000004 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111110110011,	//-0.000009 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b000000000000000000011001,	//0.000003 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b000000000000000000010100,	//0.000002 
								   24'b000000000000000000000001,	//0.000000 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b000000000000000000001111,	//0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b000000000000000000001010,	//0.000001 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b000000000000000000111000,	//0.000007 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b000000000000000000100111,	//0.000005 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b000000000000000000011111,	//0.000004 
								   24'b000000000000000000001001,	//0.000001 
								   24'b111111111111111111001100,	//-0.000006 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b000000000000000000011111,	//0.000004 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b000000000000000000100011,	//0.000004 
								   24'b000000000000000000001111,	//0.000002 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b000000000000000000001100,	//0.000001 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b000000000000000000100010,	//0.000004 
								   24'b000000000000000000000100,	//0.000000 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b000000000000000000100000,	//0.000004 
								   24'b111111111111111111001100,	//-0.000006 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b000000000000000000100110,	//0.000005 
								   24'b000000000000000000001011,	//0.000001 
								   24'b000000000000000000101000,	//0.000005 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b000000000000000000100110,	//0.000005 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111111101,	//-0.000000 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111110110110,	//-0.000009 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b000000000000000000000000,	//0.000000 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b000000000000000000010011,	//0.000002 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111011010,	//-0.000004 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b111111111111111111111010,	//-0.000001 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b000000000000000000010110,	//0.000003 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b000000000000000000000101,	//0.000001 
								   24'b111111111111111111111100,	//-0.000000 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b000000000000000000101110,	//0.000005 
								   24'b000000000000000000001000,	//0.000001 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b000000000000000000000001,	//0.000000 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111110110,	//-0.000001 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111011101,	//-0.000004 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111111000,	//-0.000001 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111011101,	//-0.000004 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111101110,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111110111,	//-0.000001 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b111111111111111111011101,	//-0.000004 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111100110,	//-0.000003 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111100000,	//-0.000004 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101011,	//-0.000002 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111111001011,	//-0.000006 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111011111,	//-0.000004 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111010011,	//-0.000005 
								   24'b111111111111111111011011,	//-0.000004 
								   24'b111111111111111111001000,	//-0.000007 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111001100,	//-0.000006 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b111111111111111111100010,	//-0.000004 
								   24'b111111111111111111101011,	//-0.000003 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111111011,	//-0.000001 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b111111111111111111110011,	//-0.000002 
								   24'b111111111111111111000011,	//-0.000007 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111001100,	//-0.000006 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111011010,	//-0.000005 
								   24'b111111111111111111101111,	//-0.000002 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111110100,	//-0.000001 
								   24'b111111111111111110111110,	//-0.000008 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111010101,	//-0.000005 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b111111111111111111010010,	//-0.000005 
								   24'b111111111111111111000110,	//-0.000007 
								   24'b111111111111111111101000,	//-0.000003 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b111111111111111111110001,	//-0.000002 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111111101010,	//-0.000003 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111010000,	//-0.000006 
								   24'b111111111111111110111011,	//-0.000008 
								   24'b111111111111111111101001,	//-0.000003 
								   24'b111111111111111110110101,	//-0.000009 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111000101,	//-0.000007 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b111111111111111111011101,	//-0.000004 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111010100,	//-0.000005 
								   24'b111111111111111111101101,	//-0.000002 
								   24'b111111111111111110110111,	//-0.000009 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b111111111111111111010111,	//-0.000005 
								   24'b111111111111111110111111,	//-0.000008 
								   24'b111111111111111111001100,	//-0.000006 
								   24'b111111111111111111000000,	//-0.000008 
								   24'b111111111111111111010001,	//-0.000006 
								   24'b111111111111111111100100,	//-0.000003 
								   24'b111111111111111111000100,	//-0.000007 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111110110001,	//-0.000009 
								   24'b111111111111111111010110,	//-0.000005 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b111111111111111111011101,	//-0.000004 
								   24'b111111111111111110110101,	//-0.000009 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111111001110,	//-0.000006 
								   24'b111111111111111111001011,	//-0.000006 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111110110001,	//-0.000009 
								   24'b111111111111111110110110,	//-0.000009 
								   24'b000000000000000000001000,	//0.000001 
								   24'b111111111111111110011101,	//-0.000012 
								   24'b111111111111111110110100,	//-0.000009 
								   24'b111111111111111111001101,	//-0.000006 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b111111111111111111011110,	//-0.000004 
								   24'b111111111111111111110011,	//-0.000001 
								   24'b111111111111111110111011,	//-0.000008 
								   24'b111111111111111111100111,	//-0.000003 
								   24'b111111111111111110110111,	//-0.000009 
								   24'b111111111111111111001010,	//-0.000006 
								   24'b111111111111111110110110,	//-0.000009 
								   24'b111111111111111111100001,	//-0.000004 
								   24'b111111111111111111000010,	//-0.000007 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111110110111,	//-0.000009 
								   24'b111111111111111110101111,	//-0.000010 
								   24'b111111111111111111000011,	//-0.000007 
								   24'b111111111111111110111001,	//-0.000008 
								   24'b111111111111111110110100,	//-0.000009 
								   24'b111111111111111110111110,	//-0.000008 
								   24'b111111111111111111000001,	//-0.000008 
								   24'b111111111111111111011000,	//-0.000005 
								   24'b111111111111111111100101,	//-0.000003 
								   24'b111111111111111110010001,	//-0.000013 
								   24'b111111111111111110000000,	//-0.000015 
								   24'b111111111111111110100101,	//-0.000011 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111110100010,	//-0.000011 
								   24'b111111111111111110110101,	//-0.000009 
								   24'b111111111111111110100000,	//-0.000011 
								   24'b111111111111111111100011,	//-0.000003 
								   24'b111111111111111111000111,	//-0.000007 
								   24'b111111111111111110010110,	//-0.000013 
								   24'b111111111111111111011001,	//-0.000005 
								   24'b111111111111111110111101,	//-0.000008 
								   24'b111111111111111111011100,	//-0.000004 
								   24'b111111111111111111111001,	//-0.000001 
								   24'b111111111111111110000101,	//-0.000015 
								   24'b111111111111111110001110,	//-0.000014 
								   24'b111111111111111110001111,	//-0.000013 
								   24'b111111111111111110010111,	//-0.000012 
								   24'b111111111111111110000100,	//-0.000015 
								   24'b111111111111111110111111,	//-0.000008 
								   24'b111111111111111110001000,	//-0.000014 
								   24'b111111111111111101111000,	//-0.000016 
								   24'b111111111111111110101000,	//-0.000011 
								   24'b111111111111111110011111,	//-0.000012 
								   24'b111111111111111110110000,	//-0.000010 
								   24'b111111111111111110010010,	//-0.000013 
								   24'b111111111111111101111110,	//-0.000016 
								   24'b111111111111111101010101,	//-0.000020 
								   24'b000000000000000000100001,	//0.000004 
								   24'b111111111111111111001111,	//-0.000006 
								   24'b111111111111111110100000,	//-0.000011 
								   24'b111111111111111101100011,	//-0.000019 
								   24'b111111111111111101010111,	//-0.000020 
								   24'b111111111111111101111100,	//-0.000016 
								   24'b000000000000000000000011,	//0.000000 
								   24'b111111111111111101111111,	//-0.000015 
								   24'b000000000000000011001110,	//0.000025 
								   24'b111111111111111101011001,	//-0.000020 
								   24'b000000000000000000000010,	//0.000000 
								   24'b111111111111111110010001,	//-0.000013 
								   24'b111111111111111110101001,	//-0.000010 
								   24'b111111111111111100111111,	//-0.000023 
								   24'b111111111111111110110001,	//-0.000009 
								   24'b000000000000000010000001,	//0.000015 
								   24'b000000000000000001010011,	//0.000010 
								   24'b111111111111111100110111,	//-0.000024 
								   24'b111111111111111110100100,	//-0.000011 
								   24'b000000000000000000000001,	//0.000000 
								   24'b000000000000000000001001,	//0.000001 
								   24'b111111111111110111101100,	//-0.000063 
								   24'b000000000000000000000110,	//0.000001 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b000000000000001000110100,	//0.000067 
								   24'b111111111111111010000000,	//-0.000046 
								   24'b111111111111111001111010,	//-0.000046 
								   24'b111111111111111011010100,	//-0.000036 
								   24'b111111111111111101100000,	//-0.000019 
								   24'b111111111111111101110001,	//-0.000017 
								   24'b111111111111111011101010,	//-0.000033 
								   24'b111111111111111100010001,	//-0.000029 
								   24'b111111111111111010111101,	//-0.000038 
								   24'b000000000000000100110101,	//0.000037 
								   24'b111111111111111111001001,	//-0.000007 
								   24'b111111111111110101000110,	//-0.000083 
								   24'b111111111111111011000010,	//-0.000038 
								   24'b111111111111110111001010,	//-0.000067 
								   24'b000000000000000111000000,	//0.000053 
								   24'b111111111111111111110000,	//-0.000002 
								   24'b111111111111111010110001,	//-0.000040 
								   24'b111111111111111110101011,	//-0.000010 
								   24'b000000000000001001011000,	//0.000072 
								   24'b111111111111111101011110,	//-0.000019 
								   24'b111111111111111111111110,	//-0.000000 
								   24'b111111111111111001100101,	//-0.000049 
								   24'b111111111111110110110001,	//-0.000070 
								   24'b111111111111101110100010,	//-0.000133 
								   24'b111111111111110100000110,	//-0.000091 
								   24'b000000000000000101100010,	//0.000042 
								   24'b000000000000000011011101,	//0.000026 
								   24'b000000000000001110101010,	//0.000112 
								   24'b111111111111111101111000,	//-0.000016 
								   24'b111111111111111011010001,	//-0.000036 
								   24'b111111111111111011010010,	//-0.000036 
								   24'b111111111111111101111011,	//-0.000016 
								   24'b000000000000000101110111,	//0.000045 
								   24'b000000000000110001011001,	//0.000377 
								   24'b111111111111111101001011,	//-0.000022 
								   24'b000000000000000111111101,	//0.000061 
								   24'b000000000000001101010100,	//0.000102 
								   24'b000000000000001111101110,	//0.000120 
								   24'b111111111111100111001000,	//-0.000190 
								   24'b111111111111110010110000,	//-0.000101 
								   24'b000000000000010001011000,	//0.000133 
								   24'b000000000000001110101110,	//0.000112 
								   24'b000000000000000101110000,	//0.000044 
								   24'b111111111111110101000111,	//-0.000083 
								   24'b111111111111111111110101,	//-0.000001 
								   24'b111111111111111011000000,	//-0.000038 
								   24'b111111111111110101010001,	//-0.000082 
								   24'b111111111111110111101010,	//-0.000064 
								   24'b111111111111111111110010,	//-0.000002 
								   24'b111111111111111000001010,	//-0.000060 
								   24'b000000000000000001110100,	//0.000014 
								   24'b000000000000001011001110,	//0.000086 
								   24'b000000000000010001001010,	//0.000131 
								   24'b000000000000010100110101,	//0.000159 
								   24'b111111111111101101001100,	//-0.000144 
								   24'b000000000000001100010101,	//0.000094 
								   24'b000000000000000001001000,	//0.000009 
								   24'b000000000000000001010010,	//0.000010 
								   24'b111111111111110011000110,	//-0.000098 
								   24'b111111111111111000001010,	//-0.000060 
								   24'b111111111111110001001000,	//-0.000113 
								   24'b000000000000000010101011,	//0.000020 
								   24'b111111111111110001010111,	//-0.000112 
								   24'b111111111111111000000001,	//-0.000061 
								   24'b111111111111111000100010,	//-0.000057 
								   24'b111111111111001100000100,	//-0.000396 
								   24'b000000000000101000011000,	//0.000308 
								   24'b000000000000001100100101,	//0.000096 
								   24'b000000000000000111011110,	//0.000057 
								   24'b000000000000001000111010,	//0.000068 
								   24'b111111111111111101011010,	//-0.000020 
								   24'b000000000000010101010100,	//0.000163 
								   24'b000000000000000000101100,	//0.000005 
								   24'b111111111111110110111110,	//-0.000069 
								   24'b000000000000010001011101,	//0.000133 
								   24'b111111111111111110101110,	//-0.000010 
								   24'b111111111111111111101100,	//-0.000002 
								   24'b000000000000001001110010,	//0.000075 
								   24'b111111111111111001000010,	//-0.000053 
								   24'b111111111111111001100110,	//-0.000049 
								   24'b000000000000011001110010,	//0.000197 
								   24'b000000000000011010000110,	//0.000199 
								   24'b111111111110111001001000,	//-0.000541 
								   24'b111111111111111011100001,	//-0.000034 
								   24'b000000000000001011000111,	//0.000085 
								   24'b000000000000000001100111,	//0.000012 
								   24'b000000000000000100010001,	//0.000033 
								   24'b111111111111110100001110,	//-0.000090 
								   24'b111111111111111011111101,	//-0.000031 
								   24'b000000000000000100101011,	//0.000036 
								   24'b000000000000011100001000,	//0.000215 
								   24'b000000000001001100010000,	//0.000582 
								   24'b111111111111110000011010,	//-0.000119 
								   24'b111111111111110101001010,	//-0.000083 
								   24'b111111111111011011011111,	//-0.000279 
								   24'b111111111111001000110011,	//-0.000421 
								   24'b111111111100101000110100,	//-0.001642 
								   24'b000000000011011000011001,	//0.001651 
								   24'b111111111100111100110000,	//-0.001490 
								   24'b000000000001000011111101,	//0.000518 
								   24'b111111111111110111110111,	//-0.000062 
								   24'b111111111111111101100001,	//-0.000019 
								   24'b111111111110111010000001,	//-0.000534 
								   24'b111111111111111110000001,	//-0.000015 
								   24'b000000000000100110010011,	//0.000292 
								   24'b000000000000001001100100,	//0.000073 
								   24'b000000000000001100100001,	//0.000096 
								   24'b111111111111111100011111,	//-0.000027 
								   24'b000000000000001010110111,	//0.000083 
								   24'b111111111111111101111110,	//-0.000015 
								   24'b111111111111111101100101,	//-0.000019 
								   24'b111111111111111110010100};	//-0.000013 
