`include "tests/eq_base_test.sv"
//`include "test/eq_simple_test.sv"
`include "tests/eq_simple_test.sv"

