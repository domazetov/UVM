//`include "sequences/eq_base_seq.sv"
`include "sequences/eq_axil_base_seq.sv"
`include "sequences/eq_axis_base_seq.sv"
//`include "sequences/eq_simple_seq.sv"
`include "sequences/eq_axil_seq.sv"
`include "sequences/eq_axis_seq.sv"

